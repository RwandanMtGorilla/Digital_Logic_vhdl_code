LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY nd2 IS
    PORT(a,b :IN STD_LOGIC;
        c :OUT STD_LOGIC);
    END;
ARCHITECTURE nd2bhv OF nd2 IS
BEGIN
    c<=a NAND b;
END;