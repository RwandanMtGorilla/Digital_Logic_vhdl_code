LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY DFF2 IS
PORT(CLK:IN STD_LOGIC;D:IN STD_LOGIC;Q:OUT STD_LOGIC);
END;
ARCHITECTURE bhv OF DFF2 IS
BEGIN
PROCESS(CLK,D)BEGIN
IF CLK='1' 
THEN Q<=D;
END IF;
END PROCESS;
END bhv;
