LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY BCD_adder1 IS
    PORT (
    BCD_A, BCD_B : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    BCD_CIN : IN STD_LOGIC;
    BCD_F : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    BCD_COUT : OUT STD_LOGIC);
END BCD_adder1;

ARCHITECTURE one OF BCD_adder1 IS
    COMPONENT full_adder_4
        PORT (
        A, B : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        F : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
        CIN : IN STD_LOGIC;
        COUT : OUT STD_LOGIC);
    END COMPONENT;

    SIGNAL temp: STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL COUT1, COUT2: STD_LOGIC;
    SIGNAL Q1, Q2: STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN
	Ul:full_adder_4 PORT MAP(A =>BCD_A,B =>BCD_B,F =>Q1,CIN =>BCD_CIN,COUT =>COUT1);
	
	COUT2<=NOT((NOT COUT1)AND(Q1(3) NAND Q1(1))AND(Q1(3)NAND Q1(2)));
	
	Q2(3)<= '0';
	Q2(2)<= COUT2;
	Q2(1)<= COUT2;
	Q2(0)<= '0';
	U2:full_adder_4 PORT MAP(A =>Q2,B =>Q1,F =>BCD_F,CIN => '0');
	
	BCD_COUT<= COUT2;
	
END one;